`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   17:28:46 04/15/2015
// Design Name:   
// Module Name:   
// Project Name:  
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: 
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module test_binary_to_grey;

	// Inputs
	reg CLK_50M;

	reg [3:0] binary;
	wire [3:0] data_out;

	binary_to_gray #(.PTR(3)) u1(
			.binary_value(binary),
			.gray_value(data_out));
	
	always
	begin
		CLK_50M=1'b0;
		#10;
		CLK_50M=1'b1;
		#10;
	end

	initial begin
		$dumpfile("grey.vcd");
		$dumpvars(data_out);
	end

	

	initial begin
		#20 binary=4'd0;
		#20 binary=4'd1;
		#20 binary=4'd2;
		#20 binary=4'd3;
		#20 binary=4'd4;
		#20 binary=4'd5;
		#20 binary=4'd6;
		#20 binary=4'd7;
		#20 binary=4'd8;
		#20 binary=4'd9;
		#20 binary=4'd10;
		#20 binary=4'd11;
		#20 binary=4'd12;
		#20 binary=4'd13;
		#20 binary=4'd14;
		#20 binary=4'd15;
		#100;$finish;
	end
      
endmodule

